* LVS netlist generated with ICnet by 'training' on Tue Dec  9 2014 at 23:18:10

*
* Globals.
*
.global GND VDD

*
* Component pathname : $MIMOS_KIT/mimos035-std-cells/schem/or02a
*
.subckt OR02A  Y A1 A0

        M4 N$431 A0 GND GND nch L=0.35u W=1.2u M=1
        M3 Y N$431 VDD VDD pch L=0.35u W=2u M=1
        M2 N$431 A1 N$429 VDD pch L=0.35u W=2u M=1
        M1 N$429 A0 VDD VDD pch L=0.35u W=2u M=1
        M6 Y N$431 GND GND nch L=0.35u W=1.2u M=1
        M5 N$431 A1 GND GND nch L=0.35u W=1.2u M=1
.ends OR02A

*
* Component pathname : $MIMOS_KIT/mimos035-std-cells/schem/and02a
*
.subckt AND02A  A1 A0 Y

        M3 Y N$647 GND GND nch L=0.35u W=1.2u M=1
        M1 N$647 A0 VDD VDD pch L=0.35u W=2u M=1
        M2 N$647 A1 VDD VDD pch L=0.35u W=2u M=1
        M4 Y N$647 VDD VDD pch L=0.35u W=2u M=1
        M5 N$647 A0 N$649 GND nch L=0.35u W=1.2u M=1
        M6 N$649 A1 GND GND nch L=0.35u W=1.2u M=1
.ends AND02A

*
* Component pathname : $MIMOS_KIT/mimos035-std-cells/schem/axor2a
*
.subckt AXOR2A  A0 A1 Y

        M9 N$470 A0 N$472 GND nch L=0.35u W=1.2u M=1
        M12 Y N$470 GND GND nch L=0.35u W=1.2u M=1
        M8 N$468 A1 GND GND nch L=0.35u W=1.2u M=1
        M7 N$467 A0 N$468 GND nch L=0.35u W=1.2u M=1
        M6 Y N$470 VDD VDD pch L=0.35u W=2u M=1
        M3 N$470 N$467 VDD VDD pch L=0.35u W=2u M=1
        M1 N$467 A0 VDD VDD pch L=0.35u W=2u M=1
        M2 N$467 A1 VDD VDD pch L=0.35u W=2u M=1
        M4 N$465 A0 VDD VDD pch L=0.35u W=2u M=1
        M5 N$470 A1 N$465 VDD pch L=0.35u W=2u M=1
        M11 N$472 N$467 GND GND nch L=0.35u W=1.2u M=1
        M10 N$470 A1 N$472 GND nch L=0.35u W=1.2u M=1
.ends AXOR2A

*
* Component pathname : /home/training/ALU_CL/schem/FullAdder
*
.subckt FULLADDER  A B COUT CIN SUM

        X_OR02A1 COUT N$21 N$18 OR02A
        X_AND02A2 CIN N$29 N$18 AND02A
        X_AND02A1 B A N$21 AND02A
        X_AXOR2A1 N$29 CIN SUM AXOR2A
        X_AXOR2A2 A B N$29 AXOR2A
.ends FULLADDER

*
* Component pathname : /home/training/ALU_CL/schem/AE
*
.subckt AE  C CIN EA A EB B WA WB AE

        X_FULLADDER1 N$38 N$40 C CIN AE FULLADDER
        X_AXOR2A3 WA N$30 N$38 AXOR2A
        X_AND02A3 A EA N$30 AND02A
        X_AXOR2A4 N$31 WB N$40 AXOR2A
        X_AND02A4 B EB N$31 AND02A
.ends AE

