* LVS netlist generated with ICnet by 'training' on Tue Dec  9 2014 at 22:01:00

*
* Globals.
*
.global GND VDD

*
* Component pathname : $MIMOS_KIT/mimos035-std-cells/schem/or02a
*
.subckt OR02A  Y A1 A0

        M4 N$431 A0 GND GND nch L=0.35u W=1.2u M=1
        M3 Y N$431 VDD VDD pch L=0.35u W=2u M=1
        M2 N$431 A1 N$429 VDD pch L=0.35u W=2u M=1
        M1 N$429 A0 VDD VDD pch L=0.35u W=2u M=1
        M6 Y N$431 GND GND nch L=0.35u W=1.2u M=1
        M5 N$431 A1 GND GND nch L=0.35u W=1.2u M=1
.ends OR02A

*
* Component pathname : $MIMOS_KIT/mimos035-std-cells/schem/and02a
*
.subckt AND02A  A1 A0 Y

        M3 Y N$647 GND GND nch L=0.35u W=1.2u M=1
        M1 N$647 A0 VDD VDD pch L=0.35u W=2u M=1
        M2 N$647 A1 VDD VDD pch L=0.35u W=2u M=1
        M4 Y N$647 VDD VDD pch L=0.35u W=2u M=1
        M5 N$647 A0 N$649 GND nch L=0.35u W=1.2u M=1
        M6 N$649 A1 GND GND nch L=0.35u W=1.2u M=1
.ends AND02A

*
* Component pathname : $MIMOS_KIT/mimos035-std-cells/schem/inv01a
*
.subckt INV01A  A Y

        M1 Y A VDD VDD pch L=0.35u W=2u M=1
        M2 Y A GND GND nch L=0.35u W=1.2u M=1
.ends INV01A

*
* Component pathname : $MIMOS_KIT/mimos035-std-cells/schem/mux21a_ni
*
.subckt MUX21A_NI  Y S0 A0 A1

        M11 N$462 A1 GND GND nch L=0.35u W=1.2u M=1
        M10 N$461 S0 N$462 GND nch L=0.35u W=1.2u M=1
        M9 N$461 N$223 N$464 GND nch L=0.35u W=1.2u M=1
        M8 Y N$461 GND GND nch L=0.35u W=1.2u M=1
        M7 N$223 S0 GND GND nch L=0.35u W=1.2u M=1
        M1 N$223 S0 VDD VDD pch L=0.35u W=2u M=1
        M4 N$459 A1 VDD VDD pch L=0.35u W=2u M=1
        M2 Y N$461 VDD VDD pch L=0.35u W=2u M=1
        M5 N$461 S0 N$457 VDD pch L=0.35u W=2u M=1
        M3 N$457 A0 VDD VDD pch L=0.35u W=2u M=1
        M12 N$464 A0 GND GND nch L=0.35u W=1.2u M=1
        M6 N$461 N$223 N$459 VDD pch L=0.35u W=2u M=1
.ends MUX21A_NI

*
* Component pathname : /home/training/ALU_CL/schem/LE
*
.subckt LE  LE S1 S2 A B

        X_OR02A1 N$21 B A OR02A
        X_AND02A1 B A N$19 AND02A
        X_INV01A1 A N$17 INV01A
        X_MUX21A_NI3 LE S2 N$10 N$9 MUX21A_NI
        X_MUX21A_NI2 N$9 S1 N$19 N$21 MUX21A_NI
        X_MUX21A_NI1 N$10 S1 A N$17 MUX21A_NI
.ends LE

