* SPICE NETLIST
***************************************

.SUBCKT MUX21a_NI S0 A0 A1 Y VDD GND
** N=28 EP=6 IP=0 FDC=12
M0 7 S0 GND GND nch L=3.5e-07 W=1.2e-06 AD=1.02e-12 AS=1.02e-12 PD=4.1e-06 PS=4.1e-06 $X=1460 $Y=3055 $D=0
M1 13 A0 GND GND nch L=3.5e-07 W=1.2e-06 AD=5.94e-13 AS=1.032e-12 PD=2.19e-06 PS=4.12e-06 $X=4130 $Y=3055 $D=0
M2 8 7 13 GND nch L=3.5e-07 W=1.2e-06 AD=6e-13 AS=5.94e-13 PD=2.2e-06 PS=2.19e-06 $X=5470 $Y=3055 $D=0
M3 14 S0 8 GND nch L=3.5e-07 W=1.2e-06 AD=5.94e-13 AS=6e-13 PD=2.19e-06 PS=2.2e-06 $X=6820 $Y=3055 $D=0
M4 GND A1 14 GND nch L=3.5e-07 W=1.2e-06 AD=1.152e-12 AS=5.94e-13 PD=4.32e-06 PS=2.19e-06 $X=8160 $Y=3055 $D=0
M5 Y 8 GND GND nch L=3.5e-07 W=1.2e-06 AD=1.02e-12 AS=1.02e-12 PD=4.1e-06 PS=4.1e-06 $X=10925 $Y=3055 $D=0
M6 7 S0 VDD VDD pch L=3.5e-07 W=2e-06 AD=1.7e-12 AS=1.7e-12 PD=5.7e-06 PS=5.7e-06 $X=1460 $Y=7925 $D=1
M7 15 A0 VDD VDD pch L=3.5e-07 W=2e-06 AD=9.75e-13 AS=1.72e-12 PD=2.975e-06 PS=5.72e-06 $X=4130 $Y=7925 $D=1
M8 8 S0 15 VDD pch L=3.5e-07 W=2e-06 AD=1.015e-12 AS=9.75e-13 PD=3.015e-06 PS=2.975e-06 $X=5455 $Y=7925 $D=1
M9 16 7 8 VDD pch L=3.5e-07 W=2e-06 AD=9.9e-13 AS=1.015e-12 PD=2.99e-06 PS=3.015e-06 $X=6820 $Y=7925 $D=1
M10 VDD A1 16 VDD pch L=3.5e-07 W=2e-06 AD=1.92e-12 AS=9.9e-13 PD=5.92e-06 PS=2.99e-06 $X=8160 $Y=7925 $D=1
M11 Y 8 VDD VDD pch L=3.5e-07 W=2e-06 AD=1.7e-12 AS=1.7e-12 PD=5.7e-06 PS=5.7e-06 $X=10925 $Y=7925 $D=1
.ENDS
***************************************
.SUBCKT LE B A S1 S2 LE VDD GND
** N=30 EP=7 IP=18 FDC=50
M0 GND 12 1 GND nch L=3.5e-07 W=1.2e-06 AD=6e-13 AS=1.2e-12 PD=2.2e-06 PS=4.4e-06 $X=-15550 $Y=1570 $D=0
M1 12 B GND GND nch L=3.5e-07 W=1.2e-06 AD=6e-13 AS=6e-13 PD=2.2e-06 PS=2.2e-06 $X=-14200 $Y=1570 $D=0
M2 GND A 12 GND nch L=3.5e-07 W=1.2e-06 AD=1.32e-12 AS=6e-13 PD=4.6e-06 PS=2.2e-06 $X=-12850 $Y=1570 $D=0
M3 GND 14 4 GND nch L=3.5e-07 W=1.2e-06 AD=6e-13 AS=1.2e-12 PD=2.2e-06 PS=4.4e-06 $X=-8040 $Y=1570 $D=0
M4 13 A GND GND nch L=3.5e-07 W=1.2e-06 AD=6e-13 AS=6e-13 PD=2.2e-06 PS=2.2e-06 $X=-6690 $Y=1570 $D=0
M5 14 B 13 GND nch L=3.5e-07 W=1.2e-06 AD=1.32e-12 AS=6e-13 PD=4.6e-06 PS=2.2e-06 $X=-5340 $Y=1570 $D=0
M6 5 A GND GND nch L=3.5e-07 W=1.2e-06 AD=1.08e-12 AS=1.02e-12 PD=4.2e-06 PS=4.1e-06 $X=-685 $Y=1570 $D=0
M7 VDD 12 1 VDD pch L=3.5e-07 W=2e-06 AD=1e-12 AS=2e-12 PD=3e-06 PS=6e-06 $X=-15550 $Y=6120 $D=1
M8 11 B VDD VDD pch L=3.5e-07 W=2e-06 AD=1e-12 AS=1e-12 PD=3e-06 PS=3e-06 $X=-14200 $Y=6120 $D=1
M9 12 A 11 VDD pch L=3.5e-07 W=2e-06 AD=2.1e-12 AS=1e-12 PD=6.1e-06 PS=3e-06 $X=-12850 $Y=6120 $D=1
M10 VDD 14 4 VDD pch L=3.5e-07 W=2e-06 AD=1e-12 AS=2e-12 PD=3e-06 PS=6e-06 $X=-8040 $Y=6120 $D=1
M11 14 A VDD VDD pch L=3.5e-07 W=2e-06 AD=1e-12 AS=1e-12 PD=3e-06 PS=3e-06 $X=-6690 $Y=6120 $D=1
M12 VDD B 14 VDD pch L=3.5e-07 W=2e-06 AD=2.1e-12 AS=1e-12 PD=6.1e-06 PS=3e-06 $X=-5340 $Y=6120 $D=1
M13 5 A VDD VDD pch L=3.5e-07 W=2e-06 AD=1.8e-12 AS=1.7e-12 PD=5.8e-06 PS=5.7e-06 $X=-685 $Y=6120 $D=1
X14 S1 A 5 8 VDD GND MUX21a_NI $T=2365 -1130 0 0 $X=1765 $Y=-3130
X15 S1 4 1 9 VDD GND MUX21a_NI $T=16295 -1130 0 0 $X=15695 $Y=-3130
X16 S2 8 9 LE VDD GND MUX21a_NI $T=30225 -1130 0 0 $X=29625 $Y=-3130
.ENDS
***************************************
