** CALIBRE LAYOUT NETLIST **
** CALIBRE VERSION: v2011.1_15.11    Thu Feb 10 17:13:25 PST 2011
** LAYOUT NAME: LE.calibre.db (LE)
** NETLIST FILE: output.spi
** GENERATED: Tue Dec  9 21:28:06 2014


.SUBCKT LE B A S1 S2 LE VDD GND 
MM0 GND 12 1 GND nch l=3.5e-07 w=1.2e-06 
MM1 12 B GND GND nch l=3.5e-07 w=1.2e-06 
MM2 GND A 12 GND nch l=3.5e-07 w=1.2e-06 
MM3 GND 14 4 GND nch l=3.5e-07 w=1.2e-06 
MM4 13 A GND GND nch l=3.5e-07 w=1.2e-06 
MM5 14 B 13 GND nch l=3.5e-07 w=1.2e-06 
MM6 5 A GND GND nch l=3.5e-07 w=1.2e-06 
MM7 VDD 12 1 VDD pch l=3.5e-07 w=2e-06 
MM8 11 B VDD VDD pch l=3.5e-07 w=2e-06 
MM9 12 A 11 VDD pch l=3.5e-07 w=2e-06 
MM10 VDD 14 4 VDD pch l=3.5e-07 w=2e-06 
MM11 14 A VDD VDD pch l=3.5e-07 w=2e-06 
MM12 VDD B 14 VDD pch l=3.5e-07 w=2e-06 
MM13 5 A VDD VDD pch l=3.5e-07 w=2e-06 
MX14/M0 X14/7 S1 GND GND nch l=3.5e-07 w=1.2e-06 
MX14/M1 X14/25 A GND GND nch l=3.5e-07 w=1.2e-06 
MX14/M2 X14/8 X14/7 X14/25 GND nch l=3.5e-07 w=1.2e-06 
MX14/M3 X14/26 S1 X14/8 GND nch l=3.5e-07 w=1.2e-06 
MX14/M4 GND 5 X14/26 GND nch l=3.5e-07 w=1.2e-06 
MX14/M5 8 X14/8 GND GND nch l=3.5e-07 w=1.2e-06 
MX14/M6 X14/7 S1 VDD VDD pch l=3.5e-07 w=2e-06 
MX14/M7 X14/27 A VDD VDD pch l=3.5e-07 w=2e-06 
MX14/M8 X14/8 S1 X14/27 VDD pch l=3.5e-07 w=2e-06 
MX14/M9 X14/28 X14/7 X14/8 VDD pch l=3.5e-07 w=2e-06 
MX14/M10 VDD 5 X14/28 VDD pch l=3.5e-07 w=2e-06 
MX14/M11 8 X14/8 VDD VDD pch l=3.5e-07 w=2e-06 
MX15/M0 X15/7 S1 GND GND nch l=3.5e-07 w=1.2e-06 
MX15/M1 X15/25 4 GND GND nch l=3.5e-07 w=1.2e-06 
MX15/M2 X15/8 X15/7 X15/25 GND nch l=3.5e-07 w=1.2e-06 
MX15/M3 X15/26 S1 X15/8 GND nch l=3.5e-07 w=1.2e-06 
MX15/M4 GND 1 X15/26 GND nch l=3.5e-07 w=1.2e-06 
MX15/M5 9 X15/8 GND GND nch l=3.5e-07 w=1.2e-06 
MX15/M6 X15/7 S1 VDD VDD pch l=3.5e-07 w=2e-06 
MX15/M7 X15/27 4 VDD VDD pch l=3.5e-07 w=2e-06 
MX15/M8 X15/8 S1 X15/27 VDD pch l=3.5e-07 w=2e-06 
MX15/M9 X15/28 X15/7 X15/8 VDD pch l=3.5e-07 w=2e-06 
MX15/M10 VDD 1 X15/28 VDD pch l=3.5e-07 w=2e-06 
MX15/M11 9 X15/8 VDD VDD pch l=3.5e-07 w=2e-06 
MX16/M0 X16/7 S2 GND GND nch l=3.5e-07 w=1.2e-06 
MX16/M1 X16/25 8 GND GND nch l=3.5e-07 w=1.2e-06 
MX16/M2 X16/8 X16/7 X16/25 GND nch l=3.5e-07 w=1.2e-06 
MX16/M3 X16/26 S2 X16/8 GND nch l=3.5e-07 w=1.2e-06 
MX16/M4 GND 9 X16/26 GND nch l=3.5e-07 w=1.2e-06 
MX16/M5 LE X16/8 GND GND nch l=3.5e-07 w=1.2e-06 
MX16/M6 X16/7 S2 VDD VDD pch l=3.5e-07 w=2e-06 
MX16/M7 X16/27 8 VDD VDD pch l=3.5e-07 w=2e-06 
MX16/M8 X16/8 S2 X16/27 VDD pch l=3.5e-07 w=2e-06 
MX16/M9 X16/28 X16/7 X16/8 VDD pch l=3.5e-07 w=2e-06 
MX16/M10 VDD 9 X16/28 VDD pch l=3.5e-07 w=2e-06 
MX16/M11 LE X16/8 VDD VDD pch l=3.5e-07 w=2e-06 
.ENDS
