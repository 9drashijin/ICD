*
* .CONNECT statements
*
.CONNECT GROUND 0
.CONNECT GND 0


* ELDO netlist generated with ICnet by 'training' on Tue Oct 14 2014 at 22:07:57

*
* Globals.
*
.global GND VDD

*
* Component pathname : $MIMOS_KIT/mimos035-std-cells/schem/axor2a
*
.subckt AXOR2A  A0 A1 Y

        M9 N$470 A0 N$472 GND nch L=0.35u W=1.2u M=1
        M12 Y N$470 GND GND nch L=0.35u W=1.2u M=1
        M8 N$468 A1 GND GND nch L=0.35u W=1.2u M=1
        M7 N$467 A0 N$468 GND nch L=0.35u W=1.2u M=1
        M6 Y N$470 VDD VDD pch L=0.35u W=2u M=1
        M3 N$470 N$467 VDD VDD pch L=0.35u W=2u M=1
        M1 N$467 A0 VDD VDD pch L=0.35u W=2u M=1
        M2 N$467 A1 VDD VDD pch L=0.35u W=2u M=1
        M4 N$465 A0 VDD VDD pch L=0.35u W=2u M=1
        M5 N$470 A1 N$465 VDD pch L=0.35u W=2u M=1
        M11 N$472 N$467 GND GND nch L=0.35u W=1.2u M=1
        M10 N$470 A1 N$472 GND nch L=0.35u W=1.2u M=1
.ends AXOR2A

*
* Component pathname : $MIMOS_KIT/mimos035-std-cells/schem/and02a
*
.subckt AND02A  A1 A0 Y

        M3 Y N$647 GND GND nch L=0.35u W=1.2u M=1
        M1 N$647 A0 VDD VDD pch L=0.35u W=2u M=1
        M2 N$647 A1 VDD VDD pch L=0.35u W=2u M=1
        M4 Y N$647 VDD VDD pch L=0.35u W=2u M=1
        M5 N$647 A0 N$649 GND nch L=0.35u W=1.2u M=1
        M6 N$649 A1 GND GND nch L=0.35u W=1.2u M=1
.ends AND02A

*
* Component pathname : $MIMOS_KIT/mimos035-std-cells/schem/or02a
*
.subckt OR02A  Y A1 A0

        M4 N$431 A0 GND GND nch L=0.35u W=1.2u M=1
        M3 Y N$431 VDD VDD pch L=0.35u W=2u M=1
        M2 N$431 A1 N$429 VDD pch L=0.35u W=2u M=1
        M1 N$429 A0 VDD VDD pch L=0.35u W=2u M=1
        M6 Y N$431 GND GND nch L=0.35u W=1.2u M=1
        M5 N$431 A1 GND GND nch L=0.35u W=1.2u M=1
.ends OR02A

*
* Component pathname : /home/training/ALU_CL/schem/FullAdder
*
.subckt FULLADDER  A B CIN COUT SUM

        X_AXOR2A2 A B N$7 AXOR2A
        X_AXOR2A1 N$7 CIN SUM AXOR2A
        X_OR02A1 COUT N$1 N$3 OR02A
        X_AND02A2 B A N$1 AND02A
        X_AND02A1 N$7 CIN N$3 AND02A
.ends FULLADDER

*
* Component pathname : /home/training/ALU_CL/schem/AE
*
.subckt AE  CIN EA A EB B WA WB AE

        X_AXOR2A2 N$1 WB N$10 AXOR2A
        X_AXOR2A1 WA N$3 N$7 AXOR2A
        X_AND02A2 B EB N$1 AND02A
        X_AND02A1 A EA N$3 AND02A
        X_FULLADDER1 N$7 N$10 CIN N$24 AE FULLADDER
.ends AE

*
* MAIN CELL: Component pathname : /home/training/ALU_CL/schem/AE_tb
*
        V8 CIN GND PULSE ( 0V 5V 1nS 1nS 1nS 60nS 120nS )
        V7 EA GND PULSE ( 0V 5V 1nS 1nS 1nS 160nS 360nS )
        V6 A GND PULSE ( 0V 5V 1nS 1nS 1nS 40nS 80nS )
        V5 EB GND PULSE ( 0V 5V 1nS 1nS 1nS 80nS 160nS )
        V4 B GND PULSE ( 0V 5V 1nS 1nS 1nS 20nS 40nS )
        V2 WB GND PULSE ( 0V 5V 1nS 1nS 1nS 20nS 40nS )
        V1 VDD GND DC 5V
        X_AE1 CIN EA A EB B GND WB AEOUT AE
*
.end
