* Component: /home/training/ALU_CL/schem/AE_tb  Viewpoint: eldonet
.INCLUDE /home/training/ALU_CL/schem/AE_tb/eldonet/AE_tb_eldonet.spi
.LIB KEY=LIB_0 $MIMOS_KIT/spice-model/035mos.eldo TYPICAL
.PROBE V




.OPTION NOASCII
.OPTION MODWL
.OPTION ENGNOT
.OPTION AEX

.TEMP 27 

.TRAN  0 1000N 0 
