*
* .CONNECT statements
*
.CONNECT GROUND 0


* ELDO netlist generated with ICnet by 'training' on Tue Nov 25 2014 at 23:16:32

*
* Globals.
*
.global VDD GND

*
* Component pathname : $MIMOS_KIT/mimos035-std-cells/schem/mux21a_ni
*
.subckt MUX21A_NI  Y S0 A0 A1

        M11 N$462 A1 GND GND nch L=0.35u W=1.2u M=1
        M10 N$461 S0 N$462 GND nch L=0.35u W=1.2u M=1
        M9 N$461 N$223 N$464 GND nch L=0.35u W=1.2u M=1
        M8 Y N$461 GND GND nch L=0.35u W=1.2u M=1
        M7 N$223 S0 GND GND nch L=0.35u W=1.2u M=1
        M1 N$223 S0 VDD VDD pch L=0.35u W=2u M=1
        M4 N$459 A1 VDD VDD pch L=0.35u W=2u M=1
        M2 Y N$461 VDD VDD pch L=0.35u W=2u M=1
        M5 N$461 S0 N$457 VDD pch L=0.35u W=2u M=1
        M3 N$457 A0 VDD VDD pch L=0.35u W=2u M=1
        M12 N$464 A0 GND GND nch L=0.35u W=1.2u M=1
        M6 N$461 N$223 N$459 VDD pch L=0.35u W=2u M=1
.ends MUX21A_NI

*
* Component pathname : $MIMOS_KIT/mimos035-std-cells/schem/and02a
*
.subckt AND02A  A1 A0 Y

        M3 Y N$647 GND GND nch L=0.35u W=1.2u M=1
        M1 N$647 A0 VDD VDD pch L=0.35u W=2u M=1
        M2 N$647 A1 VDD VDD pch L=0.35u W=2u M=1
        M4 Y N$647 VDD VDD pch L=0.35u W=2u M=1
        M5 N$647 A0 N$649 GND nch L=0.35u W=1.2u M=1
        M6 N$649 A1 GND GND nch L=0.35u W=1.2u M=1
.ends AND02A

*
* Component pathname : $MIMOS_KIT/mimos035-std-cells/schem/axor2a
*
.subckt AXOR2A  A0 A1 Y

        M9 N$470 A0 N$472 GND nch L=0.35u W=1.2u M=1
        M12 Y N$470 GND GND nch L=0.35u W=1.2u M=1
        M8 N$468 A1 GND GND nch L=0.35u W=1.2u M=1
        M7 N$467 A0 N$468 GND nch L=0.35u W=1.2u M=1
        M6 Y N$470 VDD VDD pch L=0.35u W=2u M=1
        M3 N$470 N$467 VDD VDD pch L=0.35u W=2u M=1
        M1 N$467 A0 VDD VDD pch L=0.35u W=2u M=1
        M2 N$467 A1 VDD VDD pch L=0.35u W=2u M=1
        M4 N$465 A0 VDD VDD pch L=0.35u W=2u M=1
        M5 N$470 A1 N$465 VDD pch L=0.35u W=2u M=1
        M11 N$472 N$467 GND GND nch L=0.35u W=1.2u M=1
        M10 N$470 A1 N$472 GND nch L=0.35u W=1.2u M=1
.ends AXOR2A

*
* Component pathname : /home/training/ALU_CL/schem/CE
*
.subckt CE  S0 S1 C0 S2

        X_AND02A1 S2 N$7 C0 AND02A
        X_AXOR2A1 S0 S1 N$7 AXOR2A
.ends CE

*
* Component pathname : $MIMOS_KIT/mimos035-std-cells/schem/inv01a
*
.subckt INV01A  A Y

        M1 Y A VDD VDD pch L=0.35u W=2u M=1
        M2 Y A GND GND nch L=0.35u W=1.2u M=1
.ends INV01A

*
* Component pathname : $MIMOS_KIT/mimos035-std-cells/schem/or02a
*
.subckt OR02A  Y A1 A0

        M4 N$431 A0 GND GND nch L=0.35u W=1.2u M=1
        M3 Y N$431 VDD VDD pch L=0.35u W=2u M=1
        M2 N$431 A1 N$429 VDD pch L=0.35u W=2u M=1
        M1 N$429 A0 VDD VDD pch L=0.35u W=2u M=1
        M6 Y N$431 GND GND nch L=0.35u W=1.2u M=1
        M5 N$431 A1 GND GND nch L=0.35u W=1.2u M=1
.ends OR02A

*
* Component pathname : /home/training/ALU_CL/schem/LE
*
.subckt LE  LE S1 S2 A B

        X_OR02A1 N$21 B A OR02A
        X_AND02A1 B A N$19 AND02A
        X_INV01A1 A N$17 INV01A
        X_MUX21A_NI3 LE S2 N$10 N$9 MUX21A_NI
        X_MUX21A_NI2 N$9 S1 N$19 N$21 MUX21A_NI
        X_MUX21A_NI1 N$10 S1 A N$17 MUX21A_NI
.ends LE

*
* Component pathname : /home/training/ALU_CL/schem/FullAdder
*
.subckt FULLADDER  A B CIN COUT SUM

        X_AXOR2A2 A B N$7 AXOR2A
        X_AXOR2A1 N$7 CIN SUM AXOR2A
        X_OR02A1 COUT N$1 N$3 OR02A
        X_AND02A2 B A N$1 AND02A
        X_AND02A1 N$7 CIN N$3 AND02A
.ends FULLADDER

*
* Component pathname : /home/training/ALU_CL/schem/AE
*
.subckt AE  C CIN EA A EB B WA WB AE

        X_FULLADDER1 N$38 N$40 CIN C AE FULLADDER
        X_AXOR2A3 WA N$30 N$38 AXOR2A
        X_AND02A3 A EA N$30 AND02A
        X_AXOR2A4 N$31 WB N$40 AXOR2A
        X_AND02A4 B EB N$31 AND02A
.ends AE

*
* Component pathname : /home/training/ALU_CL/schem/ALU
*
.subckt ALU  CIN COUT SUM OUT1 WB S1 S2 A B

        X_INV01A1 S1 EB INV01A
        X_MUX21A_NI1 OUT1 S2 N$3 SUM MUX21A_NI
        X_LE1 N$3 WB S1 A B LE
        X_AE1 COUT CIN VDD A EB B GND WB SUM AE
.ends ALU

*
* MAIN CELL: Component pathname : /home/training/ALU_CL/schem/ALU4bit
*
        X_MUX21A_NI2 COUT S2 N$58 N$62 MUX21A_NI
        X_MUX21A_NI1 N$62 S0 N$80 GND MUX21A_NI
        X_AND02A1 GND N$80 N$58 AND02A
        X_CE1 S0 S1 N$2 S2 CE
        X_ALU5 N$78 N$80 N$72 Q3 S0 S1 S2 A B ALU
        X_ALU7 N$2 N$99 N$103 Q0 S0 S1 S2 A B ALU
        X_ALU6 N$99 N$90 N$94 Q1 S0 S1 S2 A B ALU
        X_ALU4 N$90 N$78 N$70 Q2 S0 S1 S2 A B ALU
*
.end
