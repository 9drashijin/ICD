*
* .CONNECT statements
*
.CONNECT GROUND 0
.CONNECT GND 0


* ELDO netlist generated with ICnet by 'training' on Tue Oct 28 2014 at 21:55:07

*
* Globals.
*
.global VDD GND

*
* Component pathname : $MIMOS_KIT/mimos035-std-cells/schem/and02a
*
.subckt AND02A  A1 A0 Y

        M3 Y N$647 GND GND nch L=0.35u W=1.2u M=1
        M1 N$647 A0 VDD VDD pch L=0.35u W=2u M=1
        M2 N$647 A1 VDD VDD pch L=0.35u W=2u M=1
        M4 Y N$647 VDD VDD pch L=0.35u W=2u M=1
        M5 N$647 A0 N$649 GND nch L=0.35u W=1.2u M=1
        M6 N$649 A1 GND GND nch L=0.35u W=1.2u M=1
.ends AND02A

*
* Component pathname : $MIMOS_KIT/mimos035-std-cells/schem/axor2a
*
.subckt AXOR2A  A0 A1 Y

        M9 N$470 A0 N$472 GND nch L=0.35u W=1.2u M=1
        M12 Y N$470 GND GND nch L=0.35u W=1.2u M=1
        M8 N$468 A1 GND GND nch L=0.35u W=1.2u M=1
        M7 N$467 A0 N$468 GND nch L=0.35u W=1.2u M=1
        M6 Y N$470 VDD VDD pch L=0.35u W=2u M=1
        M3 N$470 N$467 VDD VDD pch L=0.35u W=2u M=1
        M1 N$467 A0 VDD VDD pch L=0.35u W=2u M=1
        M2 N$467 A1 VDD VDD pch L=0.35u W=2u M=1
        M4 N$465 A0 VDD VDD pch L=0.35u W=2u M=1
        M5 N$470 A1 N$465 VDD pch L=0.35u W=2u M=1
        M11 N$472 N$467 GND GND nch L=0.35u W=1.2u M=1
        M10 N$470 A1 N$472 GND nch L=0.35u W=1.2u M=1
.ends AXOR2A

*
* Component pathname : /home/training/ALU_CL/schem/CE
*
.subckt CE  S0 S1 C0 S2

        X_AND02A1 S2 N$7 C0 AND02A
        X_AXOR2A1 S0 S1 N$7 AXOR2A
.ends CE

*
* MAIN CELL: Component pathname : /home/training/ALU_CL/schem/CE_tb
*
        V4 VDD GND DC 5V
        V3 S0 GND PULSE ( 0V 5V 1nS 1nS 1nS 40nS 80nS )
        V2 S1 GND PULSE ( 0V 5V 1nS 1nS 1nS 20nS 40nS )
        V1 S2 GND PULSE ( 0V 5V 1nS 1nS 1nS 10nS 20nS )
        X_CE1 S0 S1 C0 S2 CE
*
.end
