* SPICE NETLIST
***************************************

.SUBCKT AND02a Y A0 A1 GND VDD
** N=13 EP=5 IP=0 FDC=6
M0 GND 7 Y GND nch L=3.5e-07 W=1.2e-06 AD=6e-13 AS=1.2e-12 PD=2.2e-06 PS=4.4e-06 $X=2210 $Y=2700 $D=0
M1 6 A0 GND GND nch L=3.5e-07 W=1.2e-06 AD=6e-13 AS=6e-13 PD=2.2e-06 PS=2.2e-06 $X=3560 $Y=2700 $D=0
M2 7 A1 6 GND nch L=3.5e-07 W=1.2e-06 AD=1.32e-12 AS=6e-13 PD=4.6e-06 PS=2.2e-06 $X=4910 $Y=2700 $D=0
M3 VDD 7 Y VDD pch L=3.5e-07 W=2e-06 AD=1e-12 AS=2e-12 PD=3e-06 PS=6e-06 $X=2210 $Y=7250 $D=1
M4 7 A0 VDD VDD pch L=3.5e-07 W=2e-06 AD=1e-12 AS=1e-12 PD=3e-06 PS=3e-06 $X=3560 $Y=7250 $D=1
M5 VDD A1 7 VDD pch L=3.5e-07 W=2e-06 AD=2.1e-12 AS=1e-12 PD=6.1e-06 PS=3e-06 $X=4910 $Y=7250 $D=1
.ENDS
***************************************
.SUBCKT AXOR2a A0 A1 Y GND VDD
** N=23 EP=5 IP=0 FDC=12
M0 22 A0 6 GND nch L=3.5e-07 W=1.2e-06 AD=6e-13 AS=1.2e-12 PD=2.2e-06 PS=4.4e-06 $X=1600 $Y=3100 $D=0
M1 GND A1 22 GND nch L=3.5e-07 W=1.2e-06 AD=1.2e-12 AS=6e-13 PD=4.4e-06 PS=2.2e-06 $X=2950 $Y=3100 $D=0
M2 8 A1 7 GND nch L=3.5e-07 W=1.2e-06 AD=6e-13 AS=1.2e-12 PD=2.2e-06 PS=4.4e-06 $X=5900 $Y=3000 $D=0
M3 7 A0 8 GND nch L=3.5e-07 W=1.2e-06 AD=6e-13 AS=6e-13 PD=2.2e-06 PS=2.2e-06 $X=7250 $Y=3000 $D=0
M4 GND 6 7 GND nch L=3.5e-07 W=1.2e-06 AD=1.2e-12 AS=6e-13 PD=4.4e-06 PS=2.2e-06 $X=8600 $Y=3000 $D=0
M5 Y 8 GND GND nch L=3.5e-07 W=1.2e-06 AD=1.2e-12 AS=1.2e-12 PD=4.4e-06 PS=4.4e-06 $X=11550 $Y=3000 $D=0
M6 23 A0 VDD VDD pch L=3.5e-07 W=2e-06 AD=1e-12 AS=2e-12 PD=3e-06 PS=6e-06 $X=1600 $Y=7300 $D=1
M7 8 A1 23 VDD pch L=3.5e-07 W=2e-06 AD=2e-12 AS=1e-12 PD=6e-06 PS=3e-06 $X=2950 $Y=7300 $D=1
M8 6 A1 VDD VDD pch L=3.5e-07 W=2e-06 AD=1e-12 AS=2e-12 PD=3e-06 PS=6e-06 $X=5900 $Y=7250 $D=1
M9 VDD A0 6 VDD pch L=3.5e-07 W=2e-06 AD=1e-12 AS=1e-12 PD=3e-06 PS=3e-06 $X=7250 $Y=7250 $D=1
M10 8 6 VDD VDD pch L=3.5e-07 W=2e-06 AD=2e-12 AS=1e-12 PD=6e-06 PS=3e-06 $X=8600 $Y=7250 $D=1
M11 Y 8 VDD VDD pch L=3.5e-07 W=2e-06 AD=2e-12 AS=2e-12 PD=6e-06 PS=6e-06 $X=11550 $Y=7250 $D=1
.ENDS
***************************************
.SUBCKT AE C EA A WA EB B WB CIN AE VDD GND
** N=26 EP=11 IP=40 FDC=78
M0 GND 20 C GND nch L=3.5e-07 W=1.2e-06 AD=6e-13 AS=1.2e-12 PD=2.2e-06 PS=4.4e-06 $X=52845 $Y=4735 $D=0
M1 20 2 GND GND nch L=3.5e-07 W=1.2e-06 AD=6e-13 AS=6e-13 PD=2.2e-06 PS=2.2e-06 $X=54195 $Y=4735 $D=0
M2 GND 3 20 GND nch L=3.5e-07 W=1.2e-06 AD=1.32e-12 AS=6e-13 PD=4.6e-06 PS=2.2e-06 $X=55545 $Y=4735 $D=0
M3 VDD 20 C VDD pch L=3.5e-07 W=2e-06 AD=1e-12 AS=2e-12 PD=3e-06 PS=6e-06 $X=52845 $Y=9285 $D=1
M4 19 2 VDD VDD pch L=3.5e-07 W=2e-06 AD=1e-12 AS=1e-12 PD=3e-06 PS=3e-06 $X=54195 $Y=9285 $D=1
M5 20 3 19 VDD pch L=3.5e-07 W=2e-06 AD=2.1e-12 AS=1e-12 PD=6.1e-06 PS=3e-06 $X=55545 $Y=9285 $D=1
X6 7 EA A GND VDD AND02a $T=-44770 2090 0 0 $X=-44770 $Y=90
X7 10 EB B GND VDD AND02a $T=-22555 2090 0 0 $X=-22555 $Y=90
X8 3 12 13 GND VDD AND02a $T=35615 2035 0 0 $X=35615 $Y=35
X9 2 14 CIN GND VDD AND02a $T=43130 2035 0 0 $X=43130 $Y=35
X10 WA 7 13 GND VDD AXOR2a $T=-36655 2090 0 0 $X=-37255 $Y=90
X11 10 WB 12 GND VDD AXOR2a $T=-14440 2090 0 0 $X=-15040 $Y=90
X12 12 13 14 GND VDD AXOR2a $T=6815 2035 0 0 $X=6215 $Y=35
X13 14 CIN AE GND VDD AXOR2a $T=21515 2035 0 0 $X=20915 $Y=35
.ENDS
***************************************
