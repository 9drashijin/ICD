* SPICE NETLIST
***************************************

.SUBCKT AXOR2a A0 A1 Y GND VDD
** N=23 EP=5 IP=0 FDC=12
M0 11 A0 6 GND nch L=3.5e-07 W=1.2e-06 AD=6e-13 AS=1.2e-12 PD=2.2e-06 PS=4.4e-06 $X=1600 $Y=3100 $D=0
M1 GND A1 11 GND nch L=3.5e-07 W=1.2e-06 AD=1.2e-12 AS=6e-13 PD=4.4e-06 PS=2.2e-06 $X=2950 $Y=3100 $D=0
M2 8 A1 7 GND nch L=3.5e-07 W=1.2e-06 AD=6e-13 AS=1.2e-12 PD=2.2e-06 PS=4.4e-06 $X=5900 $Y=3000 $D=0
M3 7 A0 8 GND nch L=3.5e-07 W=1.2e-06 AD=6e-13 AS=6e-13 PD=2.2e-06 PS=2.2e-06 $X=7250 $Y=3000 $D=0
M4 GND 6 7 GND nch L=3.5e-07 W=1.2e-06 AD=1.2e-12 AS=6e-13 PD=4.4e-06 PS=2.2e-06 $X=8600 $Y=3000 $D=0
M5 Y 8 GND GND nch L=3.5e-07 W=1.2e-06 AD=1.2e-12 AS=1.2e-12 PD=4.4e-06 PS=4.4e-06 $X=11550 $Y=3000 $D=0
M6 12 A0 VDD VDD pch L=3.5e-07 W=2e-06 AD=1e-12 AS=2e-12 PD=3e-06 PS=6e-06 $X=1600 $Y=7300 $D=1
M7 8 A1 12 VDD pch L=3.5e-07 W=2e-06 AD=2e-12 AS=1e-12 PD=6e-06 PS=3e-06 $X=2950 $Y=7300 $D=1
M8 6 A1 VDD VDD pch L=3.5e-07 W=2e-06 AD=1e-12 AS=2e-12 PD=3e-06 PS=6e-06 $X=5900 $Y=7250 $D=1
M9 VDD A0 6 VDD pch L=3.5e-07 W=2e-06 AD=1e-12 AS=1e-12 PD=3e-06 PS=3e-06 $X=7250 $Y=7250 $D=1
M10 8 6 VDD VDD pch L=3.5e-07 W=2e-06 AD=2e-12 AS=1e-12 PD=6e-06 PS=3e-06 $X=8600 $Y=7250 $D=1
M11 Y 8 VDD VDD pch L=3.5e-07 W=2e-06 AD=2e-12 AS=2e-12 PD=6e-06 PS=6e-06 $X=11550 $Y=7250 $D=1
.ENDS
***************************************
.SUBCKT AND02a Y A0 A1 GND VDD
** N=13 EP=5 IP=0 FDC=6
M0 GND 7 Y GND nch L=3.5e-07 W=1.2e-06 AD=6e-13 AS=1.2e-12 PD=2.2e-06 PS=4.4e-06 $X=2210 $Y=2700 $D=0
M1 6 A0 GND GND nch L=3.5e-07 W=1.2e-06 AD=6e-13 AS=6e-13 PD=2.2e-06 PS=2.2e-06 $X=3560 $Y=2700 $D=0
M2 7 A1 6 GND nch L=3.5e-07 W=1.2e-06 AD=1.32e-12 AS=6e-13 PD=4.6e-06 PS=2.2e-06 $X=4910 $Y=2700 $D=0
M3 VDD 7 Y VDD pch L=3.5e-07 W=2e-06 AD=1e-12 AS=2e-12 PD=3e-06 PS=6e-06 $X=2210 $Y=7250 $D=1
M4 7 A0 VDD VDD pch L=3.5e-07 W=2e-06 AD=1e-12 AS=1e-12 PD=3e-06 PS=3e-06 $X=3560 $Y=7250 $D=1
M5 VDD A1 7 VDD pch L=3.5e-07 W=2e-06 AD=2.1e-12 AS=1e-12 PD=6.1e-06 PS=3e-06 $X=4910 $Y=7250 $D=1
.ENDS
***************************************
.SUBCKT FullAdder COUT SUM B A CIN GND VDD
** N=18 EP=7 IP=20 FDC=42
M0 GND 10 COUT GND nch L=3.5e-07 W=1.2e-06 AD=6e-13 AS=1.2e-12 PD=2.2e-06 PS=4.4e-06 $X=28660 $Y=-490 $D=0
M1 10 2 GND GND nch L=3.5e-07 W=1.2e-06 AD=6e-13 AS=6e-13 PD=2.2e-06 PS=2.2e-06 $X=30010 $Y=-490 $D=0
M2 GND 3 10 GND nch L=3.5e-07 W=1.2e-06 AD=1.32e-12 AS=6e-13 PD=4.6e-06 PS=2.2e-06 $X=31360 $Y=-490 $D=0
M3 VDD 10 COUT VDD pch L=3.5e-07 W=2e-06 AD=1e-12 AS=2e-12 PD=3e-06 PS=6e-06 $X=28660 $Y=4060 $D=1
M4 9 2 VDD VDD pch L=3.5e-07 W=2e-06 AD=1e-12 AS=1e-12 PD=3e-06 PS=3e-06 $X=30010 $Y=4060 $D=1
M5 10 3 9 VDD pch L=3.5e-07 W=2e-06 AD=2.1e-12 AS=1e-12 PD=6.1e-06 PS=3e-06 $X=31360 $Y=4060 $D=1
X6 B A 7 GND VDD AXOR2a $T=-17370 -3190 0 0 $X=-17970 $Y=-5190
X7 7 CIN SUM GND VDD AXOR2a $T=-2670 -3190 0 0 $X=-3270 $Y=-5190
X8 3 B A GND VDD AND02a $T=11430 -3190 0 0 $X=11430 $Y=-5190
X9 2 7 CIN GND VDD AND02a $T=18945 -3190 0 0 $X=18945 $Y=-5190
.ENDS
***************************************
