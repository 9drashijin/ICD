*
* .CONNECT statements
*
.CONNECT GROUND 0
.CONNECT GND 0


* ELDO netlist generated with ICnet by 'training' on Tue Oct  7 2014 at 23:56:04

*
* Globals.
*
.global VDD GND

*
* Component pathname : $MIMOS_KIT/mimos035-std-cells/schem/axor2a
*
.subckt AXOR2A  A0 A1 Y

        M9 N$470 A0 N$472 GND nch L=0.35u W=1.2u M=1
        M12 Y N$470 GND GND nch L=0.35u W=1.2u M=1
        M8 N$468 A1 GND GND nch L=0.35u W=1.2u M=1
        M7 N$467 A0 N$468 GND nch L=0.35u W=1.2u M=1
        M6 Y N$470 VDD VDD pch L=0.35u W=2u M=1
        M3 N$470 N$467 VDD VDD pch L=0.35u W=2u M=1
        M1 N$467 A0 VDD VDD pch L=0.35u W=2u M=1
        M2 N$467 A1 VDD VDD pch L=0.35u W=2u M=1
        M4 N$465 A0 VDD VDD pch L=0.35u W=2u M=1
        M5 N$470 A1 N$465 VDD pch L=0.35u W=2u M=1
        M11 N$472 N$467 GND GND nch L=0.35u W=1.2u M=1
        M10 N$470 A1 N$472 GND nch L=0.35u W=1.2u M=1
.ends AXOR2A

*
* Component pathname : $MIMOS_KIT/mimos035-std-cells/schem/or02a
*
.subckt OR02A  Y A1 A0

        M4 N$431 A0 GND GND nch L=0.35u W=1.2u M=1
        M3 Y N$431 VDD VDD pch L=0.35u W=2u M=1
        M2 N$431 A1 N$429 VDD pch L=0.35u W=2u M=1
        M1 N$429 A0 VDD VDD pch L=0.35u W=2u M=1
        M6 Y N$431 GND GND nch L=0.35u W=1.2u M=1
        M5 N$431 A1 GND GND nch L=0.35u W=1.2u M=1
.ends OR02A

*
* Component pathname : $MIMOS_KIT/mimos035-std-cells/schem/and02a
*
.subckt AND02A  A1 A0 Y

        M3 Y N$647 GND GND nch L=0.35u W=1.2u M=1
        M1 N$647 A0 VDD VDD pch L=0.35u W=2u M=1
        M2 N$647 A1 VDD VDD pch L=0.35u W=2u M=1
        M4 Y N$647 VDD VDD pch L=0.35u W=2u M=1
        M5 N$647 A0 N$649 GND nch L=0.35u W=1.2u M=1
        M6 N$649 A1 GND GND nch L=0.35u W=1.2u M=1
.ends AND02A

*
* Component pathname : /home/training/ALU_CL/schem/FullAdder
*
.subckt FULLADDER  A B CIN COUT SUM

        X_AXOR2A2 A B N$7 AXOR2A
        X_AXOR2A1 N$7 CIN SUM AXOR2A
        X_OR02A1 COUT N$1 N$3 OR02A
        X_AND02A2 B A N$1 AND02A
        X_AND02A1 N$7 CIN N$3 AND02A
.ends FULLADDER

*
* Component pathname : /home/training/ALU_CL/schem/RippleAdder
*
.subckt RIPPLEADDER  A B S0 S1 S2 S3 COUT

        X_FULLADDER4 A B N$14 COUT S3 FULLADDER
        X_FULLADDER3 A B N$9 N$14 S2 FULLADDER
        X_FULLADDER2 A B N$38 N$9 S1 FULLADDER
        X_FULLADDER1 A B GND N$38 S0 FULLADDER
.ends RIPPLEADDER

*
* MAIN CELL: Component pathname : /home/training/ALU_CL/schem/RippleAdder_tb
*
        V3 VDD GND DC 5V
        V2 A GND PULSE ( 0V 5V 1nS 1nS 1nS 20nS 40nS )
        V1 B GND PULSE ( 0V 5V 1nS 1nS 1nS 40nS 80nS )
        X_RIPPLEADDER1 A B S0 S1 S2 S3 COUT RIPPLEADDER
*
.end
