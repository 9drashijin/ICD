* SPICE NETLIST
***************************************

.SUBCKT MUX21a_NI S0 A0 A1 Y VDD GND
** N=28 EP=6 IP=0 FDC=12
M0 7 S0 GND GND nch L=3.5e-07 W=1.2e-06 AD=1.02e-12 AS=1.02e-12 PD=4.1e-06 PS=4.1e-06 $X=1460 $Y=3055 $D=0
M1 13 A0 GND GND nch L=3.5e-07 W=1.2e-06 AD=5.94e-13 AS=1.032e-12 PD=2.19e-06 PS=4.12e-06 $X=4130 $Y=3055 $D=0
M2 8 7 13 GND nch L=3.5e-07 W=1.2e-06 AD=6e-13 AS=5.94e-13 PD=2.2e-06 PS=2.19e-06 $X=5470 $Y=3055 $D=0
M3 14 S0 8 GND nch L=3.5e-07 W=1.2e-06 AD=5.94e-13 AS=6e-13 PD=2.19e-06 PS=2.2e-06 $X=6820 $Y=3055 $D=0
M4 GND A1 14 GND nch L=3.5e-07 W=1.2e-06 AD=1.152e-12 AS=5.94e-13 PD=4.32e-06 PS=2.19e-06 $X=8160 $Y=3055 $D=0
M5 Y 8 GND GND nch L=3.5e-07 W=1.2e-06 AD=1.02e-12 AS=1.02e-12 PD=4.1e-06 PS=4.1e-06 $X=10925 $Y=3055 $D=0
M6 7 S0 VDD VDD pch L=3.5e-07 W=2e-06 AD=1.7e-12 AS=1.7e-12 PD=5.7e-06 PS=5.7e-06 $X=1460 $Y=7925 $D=1
M7 15 A0 VDD VDD pch L=3.5e-07 W=2e-06 AD=9.75e-13 AS=1.72e-12 PD=2.975e-06 PS=5.72e-06 $X=4130 $Y=7925 $D=1
M8 8 S0 15 VDD pch L=3.5e-07 W=2e-06 AD=1.015e-12 AS=9.75e-13 PD=3.015e-06 PS=2.975e-06 $X=5455 $Y=7925 $D=1
M9 16 7 8 VDD pch L=3.5e-07 W=2e-06 AD=9.9e-13 AS=1.015e-12 PD=2.99e-06 PS=3.015e-06 $X=6820 $Y=7925 $D=1
M10 VDD A1 16 VDD pch L=3.5e-07 W=2e-06 AD=1.92e-12 AS=9.9e-13 PD=5.92e-06 PS=2.99e-06 $X=8160 $Y=7925 $D=1
M11 Y 8 VDD VDD pch L=3.5e-07 W=2e-06 AD=1.7e-12 AS=1.7e-12 PD=5.7e-06 PS=5.7e-06 $X=10925 $Y=7925 $D=1
.ENDS
***************************************
.SUBCKT OR02a Y A1 A0 VDD GND
** N=13 EP=5 IP=0 FDC=6
M0 GND 7 Y GND nch L=3.5e-07 W=1.2e-06 AD=6e-13 AS=1.2e-12 PD=2.2e-06 PS=4.4e-06 $X=2100 $Y=2700 $D=0
M1 7 A1 GND GND nch L=3.5e-07 W=1.2e-06 AD=6e-13 AS=6e-13 PD=2.2e-06 PS=2.2e-06 $X=3450 $Y=2700 $D=0
M2 GND A0 7 GND nch L=3.5e-07 W=1.2e-06 AD=1.32e-12 AS=6e-13 PD=4.6e-06 PS=2.2e-06 $X=4800 $Y=2700 $D=0
M3 VDD 7 Y VDD pch L=3.5e-07 W=2e-06 AD=1e-12 AS=2e-12 PD=3e-06 PS=6e-06 $X=2100 $Y=7250 $D=1
M4 6 A1 VDD VDD pch L=3.5e-07 W=2e-06 AD=1e-12 AS=1e-12 PD=3e-06 PS=3e-06 $X=3450 $Y=7250 $D=1
M5 7 A0 6 VDD pch L=3.5e-07 W=2e-06 AD=2.1e-12 AS=1e-12 PD=6.1e-06 PS=3e-06 $X=4800 $Y=7250 $D=1
.ENDS
***************************************
.SUBCKT AND02a Y A0 A1 GND VDD
** N=13 EP=5 IP=0 FDC=6
M0 GND 7 Y GND nch L=3.5e-07 W=1.2e-06 AD=6e-13 AS=1.2e-12 PD=2.2e-06 PS=4.4e-06 $X=2210 $Y=2700 $D=0
M1 6 A0 GND GND nch L=3.5e-07 W=1.2e-06 AD=6e-13 AS=6e-13 PD=2.2e-06 PS=2.2e-06 $X=3560 $Y=2700 $D=0
M2 7 A1 6 GND nch L=3.5e-07 W=1.2e-06 AD=1.32e-12 AS=6e-13 PD=4.6e-06 PS=2.2e-06 $X=4910 $Y=2700 $D=0
M3 VDD 7 Y VDD pch L=3.5e-07 W=2e-06 AD=1e-12 AS=2e-12 PD=3e-06 PS=6e-06 $X=2210 $Y=7250 $D=1
M4 7 A0 VDD VDD pch L=3.5e-07 W=2e-06 AD=1e-12 AS=1e-12 PD=3e-06 PS=3e-06 $X=3560 $Y=7250 $D=1
M5 VDD A1 7 VDD pch L=3.5e-07 W=2e-06 AD=2.1e-12 AS=1e-12 PD=6.1e-06 PS=3e-06 $X=4910 $Y=7250 $D=1
.ENDS
***************************************
.SUBCKT AXOR2a A0 A1 Y GND VDD
** N=23 EP=5 IP=0 FDC=12
M0 11 A0 6 GND nch L=3.5e-07 W=1.2e-06 AD=6e-13 AS=1.2e-12 PD=2.2e-06 PS=4.4e-06 $X=1600 $Y=3100 $D=0
M1 GND A1 11 GND nch L=3.5e-07 W=1.2e-06 AD=1.2e-12 AS=6e-13 PD=4.4e-06 PS=2.2e-06 $X=2950 $Y=3100 $D=0
M2 8 A1 7 GND nch L=3.5e-07 W=1.2e-06 AD=6e-13 AS=1.2e-12 PD=2.2e-06 PS=4.4e-06 $X=5900 $Y=3000 $D=0
M3 7 A0 8 GND nch L=3.5e-07 W=1.2e-06 AD=6e-13 AS=6e-13 PD=2.2e-06 PS=2.2e-06 $X=7250 $Y=3000 $D=0
M4 GND 6 7 GND nch L=3.5e-07 W=1.2e-06 AD=1.2e-12 AS=6e-13 PD=4.4e-06 PS=2.2e-06 $X=8600 $Y=3000 $D=0
M5 Y 8 GND GND nch L=3.5e-07 W=1.2e-06 AD=1.2e-12 AS=1.2e-12 PD=4.4e-06 PS=4.4e-06 $X=11550 $Y=3000 $D=0
M6 12 A0 VDD VDD pch L=3.5e-07 W=2e-06 AD=1e-12 AS=2e-12 PD=3e-06 PS=6e-06 $X=1600 $Y=7300 $D=1
M7 8 A1 12 VDD pch L=3.5e-07 W=2e-06 AD=2e-12 AS=1e-12 PD=6e-06 PS=3e-06 $X=2950 $Y=7300 $D=1
M8 6 A1 VDD VDD pch L=3.5e-07 W=2e-06 AD=1e-12 AS=2e-12 PD=3e-06 PS=6e-06 $X=5900 $Y=7250 $D=1
M9 VDD A0 6 VDD pch L=3.5e-07 W=2e-06 AD=1e-12 AS=1e-12 PD=3e-06 PS=3e-06 $X=7250 $Y=7250 $D=1
M10 8 6 VDD VDD pch L=3.5e-07 W=2e-06 AD=2e-12 AS=1e-12 PD=6e-06 PS=3e-06 $X=8600 $Y=7250 $D=1
M11 Y 8 VDD VDD pch L=3.5e-07 W=2e-06 AD=2e-12 AS=2e-12 PD=6e-06 PS=6e-06 $X=11550 $Y=7250 $D=1
.ENDS
***************************************
.SUBCKT INV01a A Y VDD GND
** N=6 EP=4 IP=0 FDC=2
M0 Y A GND GND nch L=3.5e-07 W=1.2e-06 AD=1.08e-12 AS=1.02e-12 PD=4.2e-06 PS=4.1e-06 $X=2050 $Y=2700 $D=0
M1 Y A VDD VDD pch L=3.5e-07 W=2e-06 AD=1.8e-12 AS=1.7e-12 PD=5.8e-06 PS=5.7e-06 $X=2050 $Y=7250 $D=1
.ENDS
***************************************
.SUBCKT ALU VDD GND B A S1 WB CIN S2 COUT SUM OUT1
** N=25 EP=11 IP=87 FDC=142
X0 WB A 5 8 VDD GND MUX21a_NI $T=-47165 20215 0 0 $X=-47765 $Y=18215
X1 WB 6 7 9 VDD GND MUX21a_NI $T=-33235 20215 0 0 $X=-33835 $Y=18215
X2 S1 8 9 10 VDD GND MUX21a_NI $T=-19305 20215 0 0 $X=-19905 $Y=18215
X3 S2 10 SUM OUT1 VDD GND MUX21a_NI $T=109601 20215 0 0 $X=109001 $Y=18215
X4 7 B A VDD GND OR02a $T=-67180 20215 0 0 $X=-67280 $Y=18215
X5 COUT 20 21 VDD GND OR02a $T=98115 20215 0 0 $X=98015 $Y=18215
X6 6 A B GND VDD AND02a $T=-59780 20215 0 0 $X=-59780 $Y=18215
X7 12 VDD A GND VDD AND02a $T=2600 20270 0 0 $X=2600 $Y=18270
X8 14 13 B GND VDD AND02a $T=24815 20270 0 0 $X=24815 $Y=18270
X9 21 16 17 GND VDD AND02a $T=82985 20215 0 0 $X=82985 $Y=18215
X10 20 18 CIN GND VDD AND02a $T=90500 20215 0 0 $X=90500 $Y=18215
X11 GND 12 17 GND VDD AXOR2a $T=10715 20270 0 0 $X=10115 $Y=18270
X12 14 WB 16 GND VDD AXOR2a $T=32930 20270 0 0 $X=32330 $Y=18270
X13 16 17 18 GND VDD AXOR2a $T=54185 20215 0 0 $X=53585 $Y=18215
X14 18 CIN SUM GND VDD AXOR2a $T=68885 20215 0 0 $X=68285 $Y=18215
X15 A 5 VDD GND INV01a $T=-52265 20215 0 0 $X=-52265 $Y=18215
X16 S1 13 VDD GND INV01a $T=-3775 20215 0 0 $X=-3775 $Y=18215
.ENDS
***************************************
