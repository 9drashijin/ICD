** CALIBRE LAYOUT NETLIST **
** CALIBRE VERSION: v2011.1_15.11    Thu Feb 10 17:13:25 PST 2011
** LAYOUT NAME: AE.calibre.db (AE)
** NETLIST FILE: output.spi
** GENERATED: Wed Dec 10 00:35:08 2014


.SUBCKT AE C EA A WA EB B WB CIN AE VDD GND 
MM0 GND 20 C GND nch l=3.5e-07 w=1.2e-06 
MM1 20 2 GND GND nch l=3.5e-07 w=1.2e-06 
MM2 GND 3 20 GND nch l=3.5e-07 w=1.2e-06 
MM3 VDD 20 C VDD pch l=3.5e-07 w=2e-06 
MM4 19 2 VDD VDD pch l=3.5e-07 w=2e-06 
MM5 20 3 19 VDD pch l=3.5e-07 w=2e-06 
MX6/M0 GND X6/7 7 GND nch l=3.5e-07 w=1.2e-06 
MX6/M1 X6/6 EA GND GND nch l=3.5e-07 w=1.2e-06 
MX6/M2 X6/7 A X6/6 GND nch l=3.5e-07 w=1.2e-06 
MX6/M3 VDD X6/7 7 VDD pch l=3.5e-07 w=2e-06 
MX6/M4 X6/7 EA VDD VDD pch l=3.5e-07 w=2e-06 
MX6/M5 VDD A X6/7 VDD pch l=3.5e-07 w=2e-06 
MX7/M0 GND X7/7 10 GND nch l=3.5e-07 w=1.2e-06 
MX7/M1 X7/6 EB GND GND nch l=3.5e-07 w=1.2e-06 
MX7/M2 X7/7 B X7/6 GND nch l=3.5e-07 w=1.2e-06 
MX7/M3 VDD X7/7 10 VDD pch l=3.5e-07 w=2e-06 
MX7/M4 X7/7 EB VDD VDD pch l=3.5e-07 w=2e-06 
MX7/M5 VDD B X7/7 VDD pch l=3.5e-07 w=2e-06 
MX8/M0 GND X8/7 3 GND nch l=3.5e-07 w=1.2e-06 
MX8/M1 X8/6 12 GND GND nch l=3.5e-07 w=1.2e-06 
MX8/M2 X8/7 13 X8/6 GND nch l=3.5e-07 w=1.2e-06 
MX8/M3 VDD X8/7 3 VDD pch l=3.5e-07 w=2e-06 
MX8/M4 X8/7 12 VDD VDD pch l=3.5e-07 w=2e-06 
MX8/M5 VDD 13 X8/7 VDD pch l=3.5e-07 w=2e-06 
MX9/M0 GND X9/7 2 GND nch l=3.5e-07 w=1.2e-06 
MX9/M1 X9/6 14 GND GND nch l=3.5e-07 w=1.2e-06 
MX9/M2 X9/7 CIN X9/6 GND nch l=3.5e-07 w=1.2e-06 
MX9/M3 VDD X9/7 2 VDD pch l=3.5e-07 w=2e-06 
MX9/M4 X9/7 14 VDD VDD pch l=3.5e-07 w=2e-06 
MX9/M5 VDD CIN X9/7 VDD pch l=3.5e-07 w=2e-06 
MX10/M0 X10/22 WA X10/6 GND nch l=3.5e-07 w=1.2e-06 
MX10/M1 GND 7 X10/22 GND nch l=3.5e-07 w=1.2e-06 
MX10/M2 X10/8 7 X10/7 GND nch l=3.5e-07 w=1.2e-06 
MX10/M3 X10/7 WA X10/8 GND nch l=3.5e-07 w=1.2e-06 
MX10/M4 GND X10/6 X10/7 GND nch l=3.5e-07 w=1.2e-06 
MX10/M5 13 X10/8 GND GND nch l=3.5e-07 w=1.2e-06 
MX10/M6 X10/23 WA VDD VDD pch l=3.5e-07 w=2e-06 
MX10/M7 X10/8 7 X10/23 VDD pch l=3.5e-07 w=2e-06 
MX10/M8 X10/6 7 VDD VDD pch l=3.5e-07 w=2e-06 
MX10/M9 VDD WA X10/6 VDD pch l=3.5e-07 w=2e-06 
MX10/M10 X10/8 X10/6 VDD VDD pch l=3.5e-07 w=2e-06 
MX10/M11 13 X10/8 VDD VDD pch l=3.5e-07 w=2e-06 
MX11/M0 X11/22 10 X11/6 GND nch l=3.5e-07 w=1.2e-06 
MX11/M1 GND WB X11/22 GND nch l=3.5e-07 w=1.2e-06 
MX11/M2 X11/8 WB X11/7 GND nch l=3.5e-07 w=1.2e-06 
MX11/M3 X11/7 10 X11/8 GND nch l=3.5e-07 w=1.2e-06 
MX11/M4 GND X11/6 X11/7 GND nch l=3.5e-07 w=1.2e-06 
MX11/M5 12 X11/8 GND GND nch l=3.5e-07 w=1.2e-06 
MX11/M6 X11/23 10 VDD VDD pch l=3.5e-07 w=2e-06 
MX11/M7 X11/8 WB X11/23 VDD pch l=3.5e-07 w=2e-06 
MX11/M8 X11/6 WB VDD VDD pch l=3.5e-07 w=2e-06 
MX11/M9 VDD 10 X11/6 VDD pch l=3.5e-07 w=2e-06 
MX11/M10 X11/8 X11/6 VDD VDD pch l=3.5e-07 w=2e-06 
MX11/M11 12 X11/8 VDD VDD pch l=3.5e-07 w=2e-06 
MX12/M0 X12/22 12 X12/6 GND nch l=3.5e-07 w=1.2e-06 
MX12/M1 GND 13 X12/22 GND nch l=3.5e-07 w=1.2e-06 
MX12/M2 X12/8 13 X12/7 GND nch l=3.5e-07 w=1.2e-06 
MX12/M3 X12/7 12 X12/8 GND nch l=3.5e-07 w=1.2e-06 
MX12/M4 GND X12/6 X12/7 GND nch l=3.5e-07 w=1.2e-06 
MX12/M5 14 X12/8 GND GND nch l=3.5e-07 w=1.2e-06 
MX12/M6 X12/23 12 VDD VDD pch l=3.5e-07 w=2e-06 
MX12/M7 X12/8 13 X12/23 VDD pch l=3.5e-07 w=2e-06 
MX12/M8 X12/6 13 VDD VDD pch l=3.5e-07 w=2e-06 
MX12/M9 VDD 12 X12/6 VDD pch l=3.5e-07 w=2e-06 
MX12/M10 X12/8 X12/6 VDD VDD pch l=3.5e-07 w=2e-06 
MX12/M11 14 X12/8 VDD VDD pch l=3.5e-07 w=2e-06 
MX13/M0 X13/22 14 X13/6 GND nch l=3.5e-07 w=1.2e-06 
MX13/M1 GND CIN X13/22 GND nch l=3.5e-07 w=1.2e-06 
MX13/M2 X13/8 CIN X13/7 GND nch l=3.5e-07 w=1.2e-06 
MX13/M3 X13/7 14 X13/8 GND nch l=3.5e-07 w=1.2e-06 
MX13/M4 GND X13/6 X13/7 GND nch l=3.5e-07 w=1.2e-06 
MX13/M5 AE X13/8 GND GND nch l=3.5e-07 w=1.2e-06 
MX13/M6 X13/23 14 VDD VDD pch l=3.5e-07 w=2e-06 
MX13/M7 X13/8 CIN X13/23 VDD pch l=3.5e-07 w=2e-06 
MX13/M8 X13/6 CIN VDD VDD pch l=3.5e-07 w=2e-06 
MX13/M9 VDD 14 X13/6 VDD pch l=3.5e-07 w=2e-06 
MX13/M10 X13/8 X13/6 VDD VDD pch l=3.5e-07 w=2e-06 
MX13/M11 AE X13/8 VDD VDD pch l=3.5e-07 w=2e-06 
.ENDS
