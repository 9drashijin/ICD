** CALIBRE LAYOUT NETLIST **
** CALIBRE VERSION: v2011.1_15.11    Thu Feb 10 17:13:25 PST 2011
** LAYOUT NAME: ALU.calibre.db (ALU)
** NETLIST FILE: output.spi
** GENERATED: Tue Dec 16 23:05:24 2014


.SUBCKT ALU VDD GND B A S1 WB CIN S2 COUT SUM OUT1 
MX0/M0 X0/7 WB GND GND nch l=3.5e-07 w=1.2e-06 
MX0/M1 X0/25 A GND GND nch l=3.5e-07 w=1.2e-06 
MX0/M2 X0/8 X0/7 X0/25 GND nch l=3.5e-07 w=1.2e-06 
MX0/M3 X0/26 WB X0/8 GND nch l=3.5e-07 w=1.2e-06 
MX0/M4 GND 5 X0/26 GND nch l=3.5e-07 w=1.2e-06 
MX0/M5 8 X0/8 GND GND nch l=3.5e-07 w=1.2e-06 
MX0/M6 X0/7 WB VDD VDD pch l=3.5e-07 w=2e-06 
MX0/M7 X0/27 A VDD VDD pch l=3.5e-07 w=2e-06 
MX0/M8 X0/8 WB X0/27 VDD pch l=3.5e-07 w=2e-06 
MX0/M9 X0/28 X0/7 X0/8 VDD pch l=3.5e-07 w=2e-06 
MX0/M10 VDD 5 X0/28 VDD pch l=3.5e-07 w=2e-06 
MX0/M11 8 X0/8 VDD VDD pch l=3.5e-07 w=2e-06 
MX1/M0 X1/7 WB GND GND nch l=3.5e-07 w=1.2e-06 
MX1/M1 X1/25 6 GND GND nch l=3.5e-07 w=1.2e-06 
MX1/M2 X1/8 X1/7 X1/25 GND nch l=3.5e-07 w=1.2e-06 
MX1/M3 X1/26 WB X1/8 GND nch l=3.5e-07 w=1.2e-06 
MX1/M4 GND 7 X1/26 GND nch l=3.5e-07 w=1.2e-06 
MX1/M5 9 X1/8 GND GND nch l=3.5e-07 w=1.2e-06 
MX1/M6 X1/7 WB VDD VDD pch l=3.5e-07 w=2e-06 
MX1/M7 X1/27 6 VDD VDD pch l=3.5e-07 w=2e-06 
MX1/M8 X1/8 WB X1/27 VDD pch l=3.5e-07 w=2e-06 
MX1/M9 X1/28 X1/7 X1/8 VDD pch l=3.5e-07 w=2e-06 
MX1/M10 VDD 7 X1/28 VDD pch l=3.5e-07 w=2e-06 
MX1/M11 9 X1/8 VDD VDD pch l=3.5e-07 w=2e-06 
MX2/M0 X2/7 S1 GND GND nch l=3.5e-07 w=1.2e-06 
MX2/M1 X2/25 8 GND GND nch l=3.5e-07 w=1.2e-06 
MX2/M2 X2/8 X2/7 X2/25 GND nch l=3.5e-07 w=1.2e-06 
MX2/M3 X2/26 S1 X2/8 GND nch l=3.5e-07 w=1.2e-06 
MX2/M4 GND 9 X2/26 GND nch l=3.5e-07 w=1.2e-06 
MX2/M5 10 X2/8 GND GND nch l=3.5e-07 w=1.2e-06 
MX2/M6 X2/7 S1 VDD VDD pch l=3.5e-07 w=2e-06 
MX2/M7 X2/27 8 VDD VDD pch l=3.5e-07 w=2e-06 
MX2/M8 X2/8 S1 X2/27 VDD pch l=3.5e-07 w=2e-06 
MX2/M9 X2/28 X2/7 X2/8 VDD pch l=3.5e-07 w=2e-06 
MX2/M10 VDD 9 X2/28 VDD pch l=3.5e-07 w=2e-06 
MX2/M11 10 X2/8 VDD VDD pch l=3.5e-07 w=2e-06 
MX3/M0 X3/7 S2 GND GND nch l=3.5e-07 w=1.2e-06 
MX3/M1 X3/25 10 GND GND nch l=3.5e-07 w=1.2e-06 
MX3/M2 X3/8 X3/7 X3/25 GND nch l=3.5e-07 w=1.2e-06 
MX3/M3 X3/26 S2 X3/8 GND nch l=3.5e-07 w=1.2e-06 
MX3/M4 GND SUM X3/26 GND nch l=3.5e-07 w=1.2e-06 
MX3/M5 OUT1 X3/8 GND GND nch l=3.5e-07 w=1.2e-06 
MX3/M6 X3/7 S2 VDD VDD pch l=3.5e-07 w=2e-06 
MX3/M7 X3/27 10 VDD VDD pch l=3.5e-07 w=2e-06 
MX3/M8 X3/8 S2 X3/27 VDD pch l=3.5e-07 w=2e-06 
MX3/M9 X3/28 X3/7 X3/8 VDD pch l=3.5e-07 w=2e-06 
MX3/M10 VDD SUM X3/28 VDD pch l=3.5e-07 w=2e-06 
MX3/M11 OUT1 X3/8 VDD VDD pch l=3.5e-07 w=2e-06 
MX4/M0 GND X4/7 7 GND nch l=3.5e-07 w=1.2e-06 
MX4/M1 X4/7 B GND GND nch l=3.5e-07 w=1.2e-06 
MX4/M2 GND A X4/7 GND nch l=3.5e-07 w=1.2e-06 
MX4/M3 VDD X4/7 7 VDD pch l=3.5e-07 w=2e-06 
MX4/M4 X4/6 B VDD VDD pch l=3.5e-07 w=2e-06 
MX4/M5 X4/7 A X4/6 VDD pch l=3.5e-07 w=2e-06 
MX5/M0 GND X5/7 COUT GND nch l=3.5e-07 w=1.2e-06 
MX5/M1 X5/7 20 GND GND nch l=3.5e-07 w=1.2e-06 
MX5/M2 GND 21 X5/7 GND nch l=3.5e-07 w=1.2e-06 
MX5/M3 VDD X5/7 COUT VDD pch l=3.5e-07 w=2e-06 
MX5/M4 X5/6 20 VDD VDD pch l=3.5e-07 w=2e-06 
MX5/M5 X5/7 21 X5/6 VDD pch l=3.5e-07 w=2e-06 
MX6/M0 GND X6/7 6 GND nch l=3.5e-07 w=1.2e-06 
MX6/M1 X6/6 A GND GND nch l=3.5e-07 w=1.2e-06 
MX6/M2 X6/7 B X6/6 GND nch l=3.5e-07 w=1.2e-06 
MX6/M3 VDD X6/7 6 VDD pch l=3.5e-07 w=2e-06 
MX6/M4 X6/7 A VDD VDD pch l=3.5e-07 w=2e-06 
MX6/M5 VDD B X6/7 VDD pch l=3.5e-07 w=2e-06 
MX7/M0 GND X7/7 12 GND nch l=3.5e-07 w=1.2e-06 
MX7/M1 X7/6 VDD GND GND nch l=3.5e-07 w=1.2e-06 
MX7/M2 X7/7 A X7/6 GND nch l=3.5e-07 w=1.2e-06 
MX7/M3 VDD X7/7 12 VDD pch l=3.5e-07 w=2e-06 
MX7/M4 X7/7 VDD VDD VDD pch l=3.5e-07 w=2e-06 
MX7/M5 VDD A X7/7 VDD pch l=3.5e-07 w=2e-06 
MX8/M0 GND X8/7 14 GND nch l=3.5e-07 w=1.2e-06 
MX8/M1 X8/6 13 GND GND nch l=3.5e-07 w=1.2e-06 
MX8/M2 X8/7 B X8/6 GND nch l=3.5e-07 w=1.2e-06 
MX8/M3 VDD X8/7 14 VDD pch l=3.5e-07 w=2e-06 
MX8/M4 X8/7 13 VDD VDD pch l=3.5e-07 w=2e-06 
MX8/M5 VDD B X8/7 VDD pch l=3.5e-07 w=2e-06 
MX9/M0 GND X9/7 21 GND nch l=3.5e-07 w=1.2e-06 
MX9/M1 X9/6 16 GND GND nch l=3.5e-07 w=1.2e-06 
MX9/M2 X9/7 17 X9/6 GND nch l=3.5e-07 w=1.2e-06 
MX9/M3 VDD X9/7 21 VDD pch l=3.5e-07 w=2e-06 
MX9/M4 X9/7 16 VDD VDD pch l=3.5e-07 w=2e-06 
MX9/M5 VDD 17 X9/7 VDD pch l=3.5e-07 w=2e-06 
MX10/M0 GND X10/7 20 GND nch l=3.5e-07 w=1.2e-06 
MX10/M1 X10/6 18 GND GND nch l=3.5e-07 w=1.2e-06 
MX10/M2 X10/7 CIN X10/6 GND nch l=3.5e-07 w=1.2e-06 
MX10/M3 VDD X10/7 20 VDD pch l=3.5e-07 w=2e-06 
MX10/M4 X10/7 18 VDD VDD pch l=3.5e-07 w=2e-06 
MX10/M5 VDD CIN X10/7 VDD pch l=3.5e-07 w=2e-06 
MX11/M0 X11/22 GND X11/6 GND nch l=3.5e-07 w=1.2e-06 
MX11/M1 GND 12 X11/22 GND nch l=3.5e-07 w=1.2e-06 
MX11/M2 X11/8 12 X11/7 GND nch l=3.5e-07 w=1.2e-06 
MX11/M3 X11/7 GND X11/8 GND nch l=3.5e-07 w=1.2e-06 
MX11/M4 GND X11/6 X11/7 GND nch l=3.5e-07 w=1.2e-06 
MX11/M5 17 X11/8 GND GND nch l=3.5e-07 w=1.2e-06 
MX11/M6 X11/23 GND VDD VDD pch l=3.5e-07 w=2e-06 
MX11/M7 X11/8 12 X11/23 VDD pch l=3.5e-07 w=2e-06 
MX11/M8 X11/6 12 VDD VDD pch l=3.5e-07 w=2e-06 
MX11/M9 VDD GND X11/6 VDD pch l=3.5e-07 w=2e-06 
MX11/M10 X11/8 X11/6 VDD VDD pch l=3.5e-07 w=2e-06 
MX11/M11 17 X11/8 VDD VDD pch l=3.5e-07 w=2e-06 
MX12/M0 X12/22 14 X12/6 GND nch l=3.5e-07 w=1.2e-06 
MX12/M1 GND WB X12/22 GND nch l=3.5e-07 w=1.2e-06 
MX12/M2 X12/8 WB X12/7 GND nch l=3.5e-07 w=1.2e-06 
MX12/M3 X12/7 14 X12/8 GND nch l=3.5e-07 w=1.2e-06 
MX12/M4 GND X12/6 X12/7 GND nch l=3.5e-07 w=1.2e-06 
MX12/M5 16 X12/8 GND GND nch l=3.5e-07 w=1.2e-06 
MX12/M6 X12/23 14 VDD VDD pch l=3.5e-07 w=2e-06 
MX12/M7 X12/8 WB X12/23 VDD pch l=3.5e-07 w=2e-06 
MX12/M8 X12/6 WB VDD VDD pch l=3.5e-07 w=2e-06 
MX12/M9 VDD 14 X12/6 VDD pch l=3.5e-07 w=2e-06 
MX12/M10 X12/8 X12/6 VDD VDD pch l=3.5e-07 w=2e-06 
MX12/M11 16 X12/8 VDD VDD pch l=3.5e-07 w=2e-06 
MX13/M0 X13/22 16 X13/6 GND nch l=3.5e-07 w=1.2e-06 
MX13/M1 GND 17 X13/22 GND nch l=3.5e-07 w=1.2e-06 
MX13/M2 X13/8 17 X13/7 GND nch l=3.5e-07 w=1.2e-06 
MX13/M3 X13/7 16 X13/8 GND nch l=3.5e-07 w=1.2e-06 
MX13/M4 GND X13/6 X13/7 GND nch l=3.5e-07 w=1.2e-06 
MX13/M5 18 X13/8 GND GND nch l=3.5e-07 w=1.2e-06 
MX13/M6 X13/23 16 VDD VDD pch l=3.5e-07 w=2e-06 
MX13/M7 X13/8 17 X13/23 VDD pch l=3.5e-07 w=2e-06 
MX13/M8 X13/6 17 VDD VDD pch l=3.5e-07 w=2e-06 
MX13/M9 VDD 16 X13/6 VDD pch l=3.5e-07 w=2e-06 
MX13/M10 X13/8 X13/6 VDD VDD pch l=3.5e-07 w=2e-06 
MX13/M11 18 X13/8 VDD VDD pch l=3.5e-07 w=2e-06 
MX14/M0 X14/22 18 X14/6 GND nch l=3.5e-07 w=1.2e-06 
MX14/M1 GND CIN X14/22 GND nch l=3.5e-07 w=1.2e-06 
MX14/M2 X14/8 CIN X14/7 GND nch l=3.5e-07 w=1.2e-06 
MX14/M3 X14/7 18 X14/8 GND nch l=3.5e-07 w=1.2e-06 
MX14/M4 GND X14/6 X14/7 GND nch l=3.5e-07 w=1.2e-06 
MX14/M5 SUM X14/8 GND GND nch l=3.5e-07 w=1.2e-06 
MX14/M6 X14/23 18 VDD VDD pch l=3.5e-07 w=2e-06 
MX14/M7 X14/8 CIN X14/23 VDD pch l=3.5e-07 w=2e-06 
MX14/M8 X14/6 CIN VDD VDD pch l=3.5e-07 w=2e-06 
MX14/M9 VDD 18 X14/6 VDD pch l=3.5e-07 w=2e-06 
MX14/M10 X14/8 X14/6 VDD VDD pch l=3.5e-07 w=2e-06 
MX14/M11 SUM X14/8 VDD VDD pch l=3.5e-07 w=2e-06 
MX15/M0 5 A GND GND nch l=3.5e-07 w=1.2e-06 
MX15/M1 5 A VDD VDD pch l=3.5e-07 w=2e-06 
MX16/M0 13 S1 GND GND nch l=3.5e-07 w=1.2e-06 
MX16/M1 13 S1 VDD VDD pch l=3.5e-07 w=2e-06 
.ENDS
